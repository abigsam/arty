


module arty_a7_rtl (
    input  logic CLK100MHZ,
    input  logic [3:0] btn,
    input  logic [3:0] sw,
    output logic [3:0] led,
    output logic [7:0] ja
);





endmodule