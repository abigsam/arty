


module arty_a7_rtl (

);


endmodule